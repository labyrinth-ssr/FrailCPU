`include "common.svh"

module bpu(
    output i1 taken,
    input word_t resolved_branch,executed_branch,except_pc
);

    
    
endmodule