`ifndef __ADDR_TRANSLATOR
`define __ADDR_TRANSLATOR

`include "common.svh"

module addr_translator (
    input logic clk,
    input logic resetn,

    
);





endmodule

`endif
