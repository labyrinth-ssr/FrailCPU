`include "common.svh"

module pcselect(
    output word_t pc_nxt,
    input i1 branch_taken,
    input word_t pc,branch,except
);

    
    
endmodule

