`include "pipes.svh"

module pipereg2
 #(
    parameter type T=fetch_data_t
) (
    input clk,
    input reset,
    input T in[1:0],
    output T out[1:0],
    input en,flush
);
always_ff @( posedge clk ) begin
        if (reset||flush) begin 
            out[1] <= '0;
            out[0] <= '0;
        end else if (en) begin
            out <= in;
        end
    end

endmodule
