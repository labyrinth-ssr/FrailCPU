`include "Common.svh"

/**
 * NOTE: CBus does not support byte write enable mask (write_en).
 */

module DBusToCBus (
    input  dbus_req_t  dreq,
    output dbus_resp_t dresp,
    output cbus_req_t  dcreq,
    input  cbus_resp_t dcresp
);
    assign dcreq.valid    = dreq.valid;
    assign dcreq.is_write = |dreq.write_en;
    assign dcreq.order    = '0;
    assign dcreq.addr     = dreq.addr;
    assign dcreq.data     = dreq.data;

    logic okay;
    assign okay = dcresp.ready && dcresp.last;

    assign dresp.addr_ok = okay;
    assign dresp.data_ok = okay;
    assign dresp.data = dcresp.data;
endmodule
