`ifndef __MMU_SV
`define __MMU_SV

`include "common.svh"

module mmu (
    input logic clk,
    input logic resetn,

    
);





endmodule

`endif
