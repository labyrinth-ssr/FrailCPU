`include "refcpu/defs.svh"

module ExceptionReturn (
    input  context_t ctx,
    output context_t out
);
    always_comb begin
        out = ctx;
        out.state = S_FETCH;

        if (ctx.cp0.r.Status.ERL) begin
            out.pc = ctx.cp0.r.ErrorEPC;
            out.cp0.r.Status.ERL = 0;
        end else if (ctx.cp0.r.Status.EXL) begin
            out.pc = ctx.cp0.r.EPC;
            out.cp0.r.Status.EXL = 0;
        end else
            `FATAL

        if (ctx.delayed)
            `FATAL
    end
endmodule
