`ifndef __REFCPU_PKGS_SVH__
`define __REFCPU_PKGS_SVH__

`include "common.svh"

`include "refcpu/defs.svh"

`endif
